LIBRARY ieee;
--LIBRARY STD;
USE STD.textio.ALL;
USE ieee.std_logic_textio.ALL;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY SwitchTop_TB IS
END ENTITY;

ARCHITECTURE SwitchTop_TB_arc OF SwitchTop_TB IS

    COMPONENT switch_logic IS
        PORT (
            clk : IN STD_LOGIC;
            reset : IN STD_LOGIC;
            vali : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            dati : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            valo : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            dato : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;

    SIGNAL clk, reset_TB : STD_LOGIC;
    SIGNAL vali_TB, valo_TB : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL dati_TB, dato_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL COUNTER : INTEGER RANGE 0 TO 8096 := 0;
    SIGNAL PACKET1 : STD_LOGIC_VECTOR(0 TO 2247) := x"00000c9ff25794e6f7a2783f08004500010b00f44000800600000ad1f3f2174e2f54cffb005020539787ed55acd45018020046630000474554202f20485454502f312e310d0a43616368652d436f6e74726f6c3a206d61782d616765203d20333630300d0a436f6e6e656374696f6e3a204b6565702d416c6976650d0a4163636570743a202a2f2a0d0a49662d4d6f6469666965642d53696e63653a204d6f6e2c203236204a756c20323032312031363a32303a353520474d540d0a49662d4e6f6e652d4d617463683a202236306665653065372d326364220d0a557365722d4167656e743a204d6963726f736f66742d43727970746f4150492f31302e300d0a486f73743a2078312e632e6c656e63722e6f72670d0a0d0a";
    SIGNAL PACKET2 : STD_LOGIC_VECTOR(0 TO 2535) := x"94e6f7a2783f002790e6215708004500012f106140003406f002174e2f540ad1f3f20050cffbed55acd42053986a501801f5268a0000485454502f312e3120333034204e6f74204d6f6469666965640d0a436f6e74656e742d547970653a206170706c69636174696f6e2f706b69782d63726c0d0a4c6173742d4d6f6469666965643a204d6f6e2c203236204a756c20323032312031363a32303a353520474d540d0a455461673a202236306665653065372d326364220d0a43616368652d436f6e74726f6c3a206d61782d6167653d333630300d0a457870697265733a205765642c203131204d617920323032322031333a35373a343120474d540d0a446174653a205765642c203131204d617920323032322031323a35373a343120474d540d0a436f6e6e656374696f6e3a206b6565702d616c6976650d0a0d0a";
    SIGNAL PACKET3 : STD_LOGIC_VECTOR(0 TO 431) := x"00000c9ff25794e6f7a2783f08004500002800f74000800600000ad1f3f2174e2f54cffb00502053986bed55addc501001ff45800000";

BEGIN
    stimulus : PROCESS
    BEGIN
        clk <= '0';
        WAIT FOR 3 ns;
        clk <= '1';
        WAIT FOR 3 ns;
    END PROCESS;

    DUT : switch_logic PORT MAP(clk, reset_TB, vali_TB, dati_TB, valo_TB, dato_TB);

    feeder : PROCESS (clk)
    BEGIN
        IF (RISING_EDGE(clk)) THEN
            IF (COUNTER < 2240) THEN
                dati_TB(31 DOWNTO 8) <= (OTHERS => '0');
                dati_TB(7 DOWNTO 0) <= packet1(COUNTER TO COUNTER + 7);
                vali_TB(3 DOWNTO 1) <= (OTHERS => '0');
                vali_TB(0) <= '1';
                COUNTER <= COUNTER + 8;
            ELSIF (COUNTER < 2504) THEN
                dati_TB(31 DOWNTO 0) <= (OTHERS => '0');
                vali_TB(3 DOWNTO 0) <= (OTHERS => '0');
                COUNTER <= COUNTER + 8;
            ELSIF (COUNTER < 5032) THEN
                dati_TB(31 DOWNTO 16) <= (OTHERS => '0');
                dati_TB(15 DOWNTO 8) <= packet2(COUNTER - 2500 TO COUNTER - 2500 + 7);
                dati_TB(7 DOWNTO 0) <= (OTHERS => '0');
                vali_TB(3 DOWNTO 2) <= (OTHERS => '0');
                vali_TB(1) <= '1';
                vali_TB(0) <= '0';
                COUNTER <= COUNTER + 8;
            ELSIF (COUNTER < 5296) THEN
                dati_TB(31 DOWNTO 0) <= (OTHERS => '0');
                vali_TB(3 DOWNTO 0) <= (OTHERS => '0');
                COUNTER <= COUNTER + 8;
            ELSIF (COUNTER < 5728) THEN
                dati_TB(31 DOWNTO 24) <= (OTHERS => '0');
                dati_TB(23 DOWNTO 16) <= packet3(COUNTER - 5296 TO COUNTER - 5296 + 7);
                dati_TB(7 DOWNTO 0) <= (OTHERS => '0');
                vali_TB(3) <= '0';
                vali_TB(2) <= '1';
                vali_TB(1 DOWNTO 0) <= (OTHERS => '0');
                COUNTER <= COUNTER + 8;
            ELSE
                dati_TB(31 DOWNTO 0) <= (OTHERS => '0');
                vali_TB(3 DOWNTO 0) <= (OTHERS => '0');
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE;