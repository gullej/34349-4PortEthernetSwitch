LIBRARY ieee;
--LIBRARY STD;
USE STD.textio.ALL;
USE ieee.std_logic_textio.ALL;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY roundrobin_tb IS
END ENTITY;

ARCHITECTURE roundrobin_tb_arc OF roundrobin_tb IS

	COMPONENT roundrobin IS
		PORT (
			clk : IN STD_LOGIC;
			dat1 : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
			val1 : IN STD_LOGIC;
			dat2 : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
			val2 : IN STD_LOGIC;
			dat3 : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
			val3 : IN STD_LOGIC;
			dato : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			valo : OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL clk : STD_LOGIC;

	SIGNAL dat1_TB, dat2_TB, dat3_TB : STD_LOGIC_VECTOR(8 DOWNTO 0);
	SIGNAL val1_TB, val2_TB, val3_TB, valo_TB : STD_LOGIC;
	SIGNAL dato_TB : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL COUNTER : INTEGER RANGE 0 TO 1024 := 0;

	SIGNAL data1 : STD_LOGIC_VECTOR(0 TO 511) := x"180f763da5f8b831b579f47808004500028ca020400080068283c0a800b8c0265441f59e0050d9c6dba87be800c25018faf0e8280000474554202f2048545450";
	SIGNAL data2 : STD_LOGIC_VECTOR(0 TO 511) := x"2f312e310d0a486f73743a20696e736964652e6474752e646b0d0a557365722d4167656e743a204d6f7a696c6c612f352e30202857696e646f7773204e542031";
	SIGNAL data3 : STD_LOGIC_VECTOR(0 TO 511) := x"302e303b2057696e36343b207836343b2072763a39392e3029204765636b6f2f32303130303130312046697265666f782f39392e300d0a4163636570743a2074";
	SIGNAL data4 : STD_LOGIC_VECTOR(0 TO 511) := x"6578742f68746d6c2c6170706c69636174696f6e2f7868746d6c2b786d6c2c6170706c69636174696f6e2f786d6c3b713d302e392c696d6167652f617669662c";
	SIGNAL data5 : STD_LOGIC_VECTOR(0 TO 511) := x"696d6167652f776562702c2a2f2a3b713d302e380d0a4163636570742d4c616e67756167653a20656e2d55532c656e3b713d302e350d0a4163636570742d456e";
	SIGNAL data6 : STD_LOGIC_VECTOR(0 TO 511) := x"636f64696e673a20677a69702c206465666c6174650d0a444e543a20310d0a436f6e6e656374696f6e3a206b6565702d616c6976650d0a436f6f6b69653a2041";
	SIGNAL data7 : STD_LOGIC_VECTOR(0 TO 511) := x"4d43565f34443633363846343534454334313934304134433938413625343041646f62654f72673d2d323132313137393033332537434d434944545325374331";

	SIGNAL valids : STD_LOGIC_VECTOR(0 TO 63) := "0000000000000000000000000000000000000000000000000000000000000001";
BEGIN

	stimulus : PROCESS
	BEGIN
		clk <= '0';
		WAIT FOR 5 ns;
		clk <= '1';
		WAIT FOR 5 ns;
	END PROCESS;

	DUT : roundrobin PORT MAP(clk, dat1_TB, val1_TB, dat2_TB, val2_TB, dat3_TB, val3_TB, dato_TB, valo_TB);

	feeder : PROCESS (clk)
	BEGIN
		IF (RISING_EDGE(clk)) THEN
			IF (COUNTER < 64) THEN
				dat1_TB <= valids(COUNTER) & data1(COUNTER * 8 TO COUNTER * 8 + 7);
				val1_TB <= '1';
				dat2_TB <= valids(COUNTER) & data2(COUNTER * 8 TO COUNTER * 8 + 7);
				val2_TB <= '1';
				dat3_TB <= valids(COUNTER) & data3(COUNTER * 8 TO COUNTER * 8 + 7);
				val3_TB <= '1';
				COUNTER <= COUNTER + 1;
			ELSIF (COUNTER < 128) THEN
				dat1_TB <= valids(COUNTER - 64) & data4((COUNTER - 64) * 8 TO (COUNTER - 64) * 8 + 7);
				val1_TB <= '1';
				dat2_TB <= valids(COUNTER - 64) & data5((COUNTER - 64) * 8 TO (COUNTER - 64) * 8 + 7);
				val2_TB <= '1';
				dat3_TB <= valids(COUNTER - 64) & data6((COUNTER - 64) * 8 TO (COUNTER - 64) * 8 + 7);
				val3_TB <= '1';
				COUNTER <= COUNTER + 1;
			ELSIF (COUNTER < 192) THEN
				val1_TB <= '0';
				dat2_TB <= valids(COUNTER - 128) & data7((COUNTER - 128) * 8 TO (COUNTER - 128) * 8 + 7);
				val2_TB <= '1';
				val3_TB <= '0';
				COUNTER <= COUNTER + 1;
			ELSE
				val1_TB <= '0';
				val2_TB <= '0';
				val3_TB <= '0';
			END IF;
		END IF;
	END PROCESS;

END ARCHITECTURE;